//先行进位加法器
module BCLA_4 (
    ports
);
    
endmodule