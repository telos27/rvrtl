//4位比较器
module Comparator_4 (a, b, cl, ce, cg, less, equal, great);
    input [3:0] a, b;
    input cl, ce, cg;

    output less, equal, great;

    assign less = ;
    assign equal = ;
    assign great = ;
endmodule