//6到64位移位信号解码器

module ShiftDecoder_64 (datain, dataout);
    input [5:0] datain;
    output reg [63:0] dataout;

    always @(*) begin
        case(datain)
            6'b000000: dataout = 64'h0000_0000_0000_0001; 6'b000001: dataout = 64'h0000_0000_0000_0002;
            6'b000010: dataout = 64'h0000_0000_0000_0004; 6'b000011: dataout = 64'h0000_0000_0000_0008;
            6'b000100: dataout = 64'h0000_0000_0000_0010; 6'b000101: dataout = 64'h0000_0000_0000_0020;
            6'b000110: dataout = 64'h0000_0000_0000_0040; 6'b000111: dataout = 64'h0000_0000_0000_0080;
            6'b001000: dataout = 64'h0000_0000_0000_0100; 6'b001001: dataout = 64'h0000_0000_0000_0200;
            6'b001010: dataout = 64'h0000_0000_0000_0400; 6'b001011: dataout = 64'h0000_0000_0000_0800;
            6'b001100: dataout = 64'h0000_0000_0000_1000; 6'b001101: dataout = 64'h0000_0000_0000_2000;
            6'b001110: dataout = 64'h0000_0000_0000_4000; 6'b001111: dataout = 64'h0000_0000_0000_8000;
            6'b010000: dataout = 64'h0000_0000_0001_0000; 6'b010001: dataout = 64'h0000_0000_0002_0000;
            6'b010010: dataout = 64'h0000_0000_0004_0000; 6'b010011: dataout = 64'h0000_0000_0008_0000;
            6'b010100: dataout = 64'h0000_0000_0010_0000; 6'b010101: dataout = 64'h0000_0000_0020_0000;
            6'b010110: dataout = 64'h0000_0000_0040_0000; 6'b010111: dataout = 64'h0000_0000_0080_0000;
            6'b011000: dataout = 64'h0000_0000_0100_0000; 6'b011001: dataout = 64'h0000_0000_0200_0000;
            6'b011010: dataout = 64'h0000_0000_0400_0000; 6'b011011: dataout = 64'h0000_0000_0800_0000;
            6'b011100: dataout = 64'h0000_0000_1000_0000; 6'b011101: dataout = 64'h0000_0000_2000_0000;
            6'b011110: dataout = 64'h0000_0000_4000_0000; 6'b011111: dataout = 64'h0000_0000_8000_0000;
            6'b100000: dataout = 64'h0000_0001_0000_0000; 6'b100001: dataout = 64'h0000_0002_0000_0000;
            6'b100010: dataout = 64'h0000_0004_0000_0000; 6'b100011: dataout = 64'h0000_0008_0000_0000;
            6'b100100: dataout = 64'h0000_0010_0000_0000; 6'b100101: dataout = 64'h0000_0020_0000_0000;
            6'b100110: dataout = 64'h0000_0040_0000_0000; 6'b100111: dataout = 64'h0000_0080_0000_0000;
            6'b101000: dataout = 64'h0000_0100_0000_0000; 6'b101001: dataout = 64'h0000_0200_0000_0000;
            6'b101010: dataout = 64'h0000_0400_0000_0000; 6'b101011: dataout = 64'h0000_0800_0000_0000;
            6'b101100: dataout = 64'h0000_1000_0000_0000; 6'b101101: dataout = 64'h0000_2000_0000_0000;
            6'b101110: dataout = 64'h0000_4000_0000_0000; 6'b101111: dataout = 64'h0000_8000_0000_0000;
            6'b110000: dataout = 64'h0001_0000_0000_0000; 6'b110001: dataout = 64'h0002_0000_0000_0000;
            6'b110010: dataout = 64'h0004_0000_0000_0000; 6'b110011: dataout = 64'h0008_0000_0000_0000;
            6'b110100: dataout = 64'h0010_0000_0000_0000; 6'b110101: dataout = 64'h0020_0000_0000_0000;
            6'b110110: dataout = 64'h0040_0000_0000_0000; 6'b110111: dataout = 64'h0080_0000_0000_0000;
            6'b111000: dataout = 64'h0100_0000_0000_0000; 6'b111001: dataout = 64'h0200_0000_0000_0000;
            6'b111010: dataout = 64'h0400_0000_0000_0000; 6'b111011: dataout = 64'h0800_0000_0000_0000;
            6'b111100: dataout = 64'h1000_0000_0000_0000; 6'b111101: dataout = 64'h2000_0000_0000_0000;
            6'b111110: dataout = 64'h4000_0000_0000_0000; 6'b111111: dataout = 64'h8000_0000_0000_0000;
            default: dataout = 64'h0000_0000_0000_0000;
        endcase
    end

endmodule