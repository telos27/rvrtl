//移位信号生成
module Shift_Signal (shift5, shift32);
    input [4:0] shift5;
    output reg [31:0] shift32;

    always @(*) begin
    case (s)
        //0~3
        5'b00000: shift = 32'h0000_0001;
        5'b00001: shift = 32'h0000_0002;
        5'b00010: shift = 32'h0000_0004;
        5'b00011: shift = 32'h0000_0008;
        //4~7
        5'b00100: shift = 32'h0000_0010;
        5'b00101: shift = 32'h0000_0020;
        5'b00110: shift = 32'h0000_0040;
        5'b00111: shift = 32'h0000_0080;
        //8~11
        5'b01000: shift = 32'h0000_0100;
        5'b01001: shift = 32'h0000_0200;
        5'b01010: shift = 32'h0000_0400;
        5'b01011: shift = 32'h0000_0800;
        //12~15
        5'b01100: shift = 32'h0000_1000;
        5'b01101: shift = 32'h0000_2000;
        5'b01110: shift = 32'h0000_4000;
        5'b01111: shift = 32'h0000_8000;
        //16~19
        5'b10000: shift = 32'h0001_0000;
        5'b10001: shift = 32'h0002_0000;
        5'b10010: shift = 32'h0004_0000;
        5'b10011: shift = 32'h0008_0000;
        //20~23
        5'b10100: shift = 32'h0010_0000;
        5'b10101: shift = 32'h0020_0000;
        5'b10110: shift = 32'h0040_0000;
        5'b10111: shift = 32'h0080_0000;
        //24~27
        5'b11000: shift = 32'h0100_0000;
        5'b11001: shift = 32'h0200_0000;
        5'b11010: shift = 32'h0400_0000;
        5'b11011: shift = 32'h0800_0000;
        //28~31
        5'b11100: shift = 32'h1000_0000;
        5'b11101: shift = 32'h2000_0000;
        5'b11110: shift = 32'h4000_0000;
        5'b11111: shift = 32'h8000_0000;
    endcase
    end
endmodule
